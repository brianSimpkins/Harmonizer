module fft(input logic sck, sdi,
			  output logic sdo, done);
			  
	// Create spi module, input module, output module
	
	// Route SPI buffer to FFT input
	
	// Route FFT output to SPI buffer
	
	// Have logic which waits until SPI is full before starting FFT inputting
	
	// Have logic which, once FFT output is full, pulses reset in the FFT
	
endmodule