module spi();
endmodule